*test_mos devices

m0 vdn vgn 0 vbn NMOS_VTL L=45e-9 W=360e-9
m1 0 vgp vdp vbp PMOS_VTL L=45e-9 W=360e-9
.END
