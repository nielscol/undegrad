* SPICE NETLIST
***************************************

.SUBCKT adder A_15 A_14 A_13 A_12 A_11 A_10 A_9 A_8 A_7 A_6 A_5 A_4 A_3 A_2 A_1 A_0 B_15 B_14 B_13 B_12
+ B_11 B_10 B_9 B_8 B_7 B_6 B_5 B_4 B_3 B_2 B_1 B_0 GND! S_0 Cout VDD! S_15 S_14 S_13 S_12
+ S_11 S_10 S_9 S_8 S_7 S_6 S_5 S_4 S_3 S_2 S_1
** N=476 EP=51 IP=0 FDC=884
M0 119 A_15 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=-8250 $D=1
M1 380 A_15 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=-3800 $D=1
M2 121 A_14 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=650 $D=1
M3 381 A_14 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=5100 $D=1
M4 123 A_13 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=9550 $D=1
M5 382 A_13 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=14000 $D=1
M6 125 A_12 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=18450 $D=1
M7 383 A_12 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=22900 $D=1
M8 127 A_11 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=27350 $D=1
M9 384 A_11 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=31800 $D=1
M10 129 A_10 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=36250 $D=1
M11 385 A_10 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=40700 $D=1
M12 131 A_9 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=45150 $D=1
M13 386 A_9 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=49600 $D=1
M14 133 A_8 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=54050 $D=1
M15 387 A_8 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=58500 $D=1
M16 135 A_7 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=62950 $D=1
M17 388 A_7 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=67400 $D=1
M18 137 A_6 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=71850 $D=1
M19 389 A_6 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=76300 $D=1
M20 139 A_5 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=80750 $D=1
M21 390 A_5 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=85200 $D=1
M22 141 A_4 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=89650 $D=1
M23 391 A_4 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=94100 $D=1
M24 143 A_3 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=98550 $D=1
M25 392 A_3 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=103000 $D=1
M26 145 A_2 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=107450 $D=1
M27 393 A_2 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=111900 $D=1
M28 147 A_1 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=116350 $D=1
M29 394 A_1 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=120800 $D=1
M30 149 A_0 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=125250 $D=1
M31 395 A_0 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=450 $Y=129700 $D=1
M32 GND! B_15 119 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=-8250 $D=1
M33 120 B_15 380 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=-3800 $D=1
M34 GND! B_14 121 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=650 $D=1
M35 122 B_14 381 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=5100 $D=1
M36 GND! B_13 123 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=9550 $D=1
M37 124 B_13 382 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=14000 $D=1
M38 GND! B_12 125 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=18450 $D=1
M39 126 B_12 383 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=22900 $D=1
M40 GND! B_11 127 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=27350 $D=1
M41 128 B_11 384 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=31800 $D=1
M42 GND! B_10 129 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=36250 $D=1
M43 130 B_10 385 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=40700 $D=1
M44 GND! B_9 131 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=45150 $D=1
M45 132 B_9 386 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=49600 $D=1
M46 GND! B_8 133 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=54050 $D=1
M47 134 B_8 387 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=58500 $D=1
M48 GND! B_7 135 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=62950 $D=1
M49 136 B_7 388 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=67400 $D=1
M50 GND! B_6 137 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=71850 $D=1
M51 138 B_6 389 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=76300 $D=1
M52 GND! B_5 139 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=80750 $D=1
M53 140 B_5 390 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=85200 $D=1
M54 GND! B_4 141 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=89650 $D=1
M55 142 B_4 391 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=94100 $D=1
M56 GND! B_3 143 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=98550 $D=1
M57 144 B_3 392 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=103000 $D=1
M58 GND! B_2 145 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=107450 $D=1
M59 146 B_2 393 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=111900 $D=1
M60 GND! B_1 147 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=116350 $D=1
M61 148 B_1 394 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=120800 $D=1
M62 GND! B_0 149 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=125250 $D=1
M63 150 B_0 395 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=900 $Y=129700 $D=1
M64 GND! 119 41 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=-8250 $D=1
M65 GND! 121 33 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=650 $D=1
M66 GND! 123 34 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=9550 $D=1
M67 GND! 125 35 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=18450 $D=1
M68 GND! 127 42 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=27350 $D=1
M69 GND! 129 36 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=36250 $D=1
M70 GND! 131 43 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=45150 $D=1
M71 GND! 133 37 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=54050 $D=1
M72 GND! 135 44 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=62950 $D=1
M73 GND! 137 38 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=71850 $D=1
M74 GND! 139 45 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=80750 $D=1
M75 GND! 141 39 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=89650 $D=1
M76 GND! 143 46 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=98550 $D=1
M77 GND! 145 40 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=107450 $D=1
M78 GND! 147 47 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=116350 $D=1
M79 GND! 149 55 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=1800 $Y=125250 $D=1
M80 151 120 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=-3800 $D=1
M81 152 122 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=5100 $D=1
M82 48 124 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=14000 $D=1
M83 153 126 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=22900 $D=1
M84 49 128 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=31800 $D=1
M85 154 130 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=40700 $D=1
M86 50 132 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=49600 $D=1
M87 155 134 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=58500 $D=1
M88 51 136 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=67400 $D=1
M89 156 138 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=76300 $D=1
M90 52 140 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=85200 $D=1
M91 157 142 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=94100 $D=1
M92 53 144 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=103000 $D=1
M93 158 146 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=111900 $D=1
M94 54 148 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=120800 $D=1
M95 159 150 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1900 $Y=129700 $D=1
M96 396 A_15 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=-8250 $D=1
M97 397 A_14 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=650 $D=1
M98 398 A_13 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=9550 $D=1
M99 399 A_12 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=18450 $D=1
M100 400 A_11 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=27350 $D=1
M101 401 A_10 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=36250 $D=1
M102 402 A_9 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=45150 $D=1
M103 403 A_8 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=54050 $D=1
M104 404 A_7 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=62950 $D=1
M105 405 A_6 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=71850 $D=1
M106 406 A_5 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=80750 $D=1
M107 407 A_4 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=89650 $D=1
M108 408 A_3 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=98550 $D=1
M109 409 A_2 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=107450 $D=1
M110 410 A_1 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=116350 $D=1
M111 411 A_0 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=2250 $Y=125250 $D=1
M112 41 B_15 396 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=-8250 $D=1
M113 33 B_14 397 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=650 $D=1
M114 34 B_13 398 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=9550 $D=1
M115 35 B_12 399 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=18450 $D=1
M116 42 B_11 400 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=27350 $D=1
M117 36 B_10 401 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=36250 $D=1
M118 43 B_9 402 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=45150 $D=1
M119 37 B_8 403 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=54050 $D=1
M120 44 B_7 404 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=62950 $D=1
M121 38 B_6 405 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=71850 $D=1
M122 45 B_5 406 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=80750 $D=1
M123 39 B_4 407 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=89650 $D=1
M124 46 B_3 408 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=98550 $D=1
M125 40 B_2 409 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=107450 $D=1
M126 47 B_1 410 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=116350 $D=1
M127 55 B_0 411 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=2700 $Y=125250 $D=1
M128 412 34 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=650 $D=1
M129 176 152 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=5100 $D=1
M130 177 34 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=9550 $D=1
M131 178 48 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=14000 $D=1
M132 413 42 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=18450 $D=1
M133 179 153 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=22900 $D=1
M134 180 42 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=27350 $D=1
M135 181 49 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=31800 $D=1
M136 414 43 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=36250 $D=1
M137 182 154 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=40700 $D=1
M138 183 43 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=45150 $D=1
M139 184 50 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=49600 $D=1
M140 415 44 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=54050 $D=1
M141 185 155 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=58500 $D=1
M142 186 44 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=62950 $D=1
M143 187 51 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=67400 $D=1
M144 416 45 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=71850 $D=1
M145 188 156 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=76300 $D=1
M146 189 45 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=80750 $D=1
M147 190 52 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=85200 $D=1
M148 417 46 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=89650 $D=1
M149 191 157 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=94100 $D=1
M150 192 46 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=98550 $D=1
M151 193 53 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=103000 $D=1
M152 418 47 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=107450 $D=1
M153 194 158 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=111900 $D=1
M154 195 47 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=116350 $D=1
M155 196 54 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=3700 $Y=120800 $D=1
M156 197 159 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=3700 $Y=129700 $D=1
M157 198 33 412 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=4150 $Y=650 $D=1
M158 419 33 176 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=4150 $Y=5100 $D=1
M159 199 35 413 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=4150 $Y=18450 $D=1
M160 420 35 179 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=4150 $Y=22900 $D=1
M161 200 36 414 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=4150 $Y=36250 $D=1
M162 421 36 182 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=4150 $Y=40700 $D=1
M163 201 37 415 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=4150 $Y=54050 $D=1
M164 422 37 185 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=4150 $Y=58500 $D=1
M165 202 38 416 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=4150 $Y=71850 $D=1
M166 423 38 188 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=4150 $Y=76300 $D=1
M167 203 39 417 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=4150 $Y=89650 $D=1
M168 424 39 191 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=4150 $Y=94100 $D=1
M169 204 40 418 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=4150 $Y=107450 $D=1
M170 425 40 194 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=4150 $Y=111900 $D=1
M171 426 55 197 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=4150 $Y=129700 $D=1
M172 GND! 48 419 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=4600 $Y=5100 $D=1
M173 GND! 49 420 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=4600 $Y=22900 $D=1
M174 GND! 50 421 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=4600 $Y=40700 $D=1
M175 GND! 51 422 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=4600 $Y=58500 $D=1
M176 GND! 52 423 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=4600 $Y=76300 $D=1
M177 GND! 53 424 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=4600 $Y=94100 $D=1
M178 GND! 54 425 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=4600 $Y=111900 $D=1
M179 GND! GND! 426 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=4600 $Y=129700 $D=1
M180 57 177 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=9550 $D=1
M181 213 178 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=14000 $D=1
M182 58 180 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=27350 $D=1
M183 214 181 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=31800 $D=1
M184 59 183 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=45150 $D=1
M185 215 184 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=49600 $D=1
M186 60 186 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=62950 $D=1
M187 216 187 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=67400 $D=1
M188 61 189 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=80750 $D=1
M189 217 190 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=85200 $D=1
M190 62 192 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=98550 $D=1
M191 218 193 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=103000 $D=1
M192 63 195 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=116350 $D=1
M193 219 196 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=4700 $Y=120800 $D=1
M194 64 198 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=5150 $Y=650 $D=1
M195 65 199 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=5150 $Y=18450 $D=1
M196 66 200 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=5150 $Y=36250 $D=1
M197 67 201 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=5150 $Y=54050 $D=1
M198 68 202 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=5150 $Y=71850 $D=1
M199 69 203 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=5150 $Y=89650 $D=1
M200 70 204 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=5150 $Y=107450 $D=1
M201 220 176 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=5500 $Y=5100 $D=1
M202 71 179 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=5500 $Y=22900 $D=1
M203 72 182 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=5500 $Y=40700 $D=1
M204 73 185 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=5500 $Y=58500 $D=1
M205 74 188 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=5500 $Y=76300 $D=1
M206 75 191 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=5500 $Y=94100 $D=1
M207 76 194 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=5500 $Y=111900 $D=1
M208 77 197 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=5500 $Y=129700 $D=1
M209 427 65 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=650 $D=1
M210 221 220 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=5100 $D=1
M211 428 66 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=18450 $D=1
M212 222 71 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=22900 $D=1
M213 429 67 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=36250 $D=1
M214 223 72 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=40700 $D=1
M215 430 68 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=54050 $D=1
M216 224 73 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=58500 $D=1
M217 431 69 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=71850 $D=1
M218 225 74 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=76300 $D=1
M219 432 70 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=89650 $D=1
M220 226 75 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=94100 $D=1
M221 227 76 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=6500 $Y=111900 $D=1
M222 228 55 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=6500 $Y=125250 $D=1
M223 229 77 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=6500 $Y=129700 $D=1
M224 230 64 427 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=6950 $Y=650 $D=1
M225 433 64 221 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=6950 $Y=5100 $D=1
M226 231 65 428 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=6950 $Y=18450 $D=1
M227 434 65 222 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=6950 $Y=22900 $D=1
M228 232 66 429 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=6950 $Y=36250 $D=1
M229 435 66 223 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=6950 $Y=40700 $D=1
M230 233 67 430 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=6950 $Y=54050 $D=1
M231 436 67 224 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=6950 $Y=58500 $D=1
M232 234 68 431 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=6950 $Y=71850 $D=1
M233 437 68 225 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=6950 $Y=76300 $D=1
M234 235 69 432 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=6950 $Y=89650 $D=1
M235 438 69 226 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=6950 $Y=94100 $D=1
M236 439 70 227 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=6950 $Y=111900 $D=1
M237 GND! 71 433 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=7400 $Y=5100 $D=1
M238 GND! 72 434 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=7400 $Y=22900 $D=1
M239 GND! 73 435 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=7400 $Y=40700 $D=1
M240 GND! 74 436 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=7400 $Y=58500 $D=1
M241 GND! 75 437 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=7400 $Y=76300 $D=1
M242 GND! 76 438 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=7400 $Y=94100 $D=1
M243 GND! 77 439 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=7400 $Y=111900 $D=1
M244 S_0 228 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=7500 $Y=125250 $D=1
M245 89 229 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=7500 $Y=129700 $D=1
M246 78 230 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=7950 $Y=650 $D=1
M247 79 231 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=7950 $Y=18450 $D=1
M248 80 232 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=7950 $Y=36250 $D=1
M249 81 233 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=7950 $Y=54050 $D=1
M250 82 234 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=7950 $Y=71850 $D=1
M251 83 235 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=7950 $Y=89650 $D=1
M252 244 221 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=8300 $Y=5100 $D=1
M253 245 222 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=8300 $Y=22900 $D=1
M254 87 223 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=8300 $Y=40700 $D=1
M255 85 224 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=8300 $Y=58500 $D=1
M256 84 225 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=8300 $Y=76300 $D=1
M257 88 226 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=8300 $Y=94100 $D=1
M258 86 227 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=8300 $Y=111900 $D=1
M259 440 80 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=650 $D=1
M260 246 244 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=5100 $D=1
M261 441 81 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=18450 $D=1
M262 247 245 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=22900 $D=1
M263 442 82 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=36250 $D=1
M264 248 87 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=40700 $D=1
M265 443 83 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=54050 $D=1
M266 249 85 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=58500 $D=1
M267 250 84 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=76300 $D=1
M268 251 88 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=9300 $Y=94100 $D=1
M269 252 40 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=9300 $Y=107450 $D=1
M270 253 86 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=9300 $Y=111900 $D=1
M271 254 78 440 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=9750 $Y=650 $D=1
M272 444 78 246 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=9750 $Y=5100 $D=1
M273 255 79 441 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=9750 $Y=18450 $D=1
M274 445 79 247 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=9750 $Y=22900 $D=1
M275 256 80 442 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=9750 $Y=36250 $D=1
M276 446 80 248 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=9750 $Y=40700 $D=1
M277 257 81 443 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=9750 $Y=54050 $D=1
M278 447 81 249 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=9750 $Y=58500 $D=1
M279 448 82 250 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=9750 $Y=76300 $D=1
M280 449 83 251 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=9750 $Y=94100 $D=1
M281 GND! 87 444 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=10200 $Y=5100 $D=1
M282 GND! 85 445 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=10200 $Y=22900 $D=1
M283 GND! 84 446 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=10200 $Y=40700 $D=1
M284 GND! 88 447 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=10200 $Y=58500 $D=1
M285 GND! 86 448 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=10200 $Y=76300 $D=1
M286 GND! 89 449 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=10200 $Y=94100 $D=1
M287 107 252 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=10300 $Y=107450 $D=1
M288 96 253 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=10300 $Y=111900 $D=1
M289 90 254 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=10750 $Y=650 $D=1
M290 91 255 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=10750 $Y=18450 $D=1
M291 92 256 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=10750 $Y=36250 $D=1
M292 93 257 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=10750 $Y=54050 $D=1
M293 264 246 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=11100 $Y=5100 $D=1
M294 265 247 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=11100 $Y=22900 $D=1
M295 266 248 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=11100 $Y=40700 $D=1
M296 267 249 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=11100 $Y=58500 $D=1
M297 94 250 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=11100 $Y=76300 $D=1
M298 95 251 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=11100 $Y=94100 $D=1
M299 268 264 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=12100 $Y=5100 $D=1
M300 269 265 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=12100 $Y=22900 $D=1
M301 270 266 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=12100 $Y=40700 $D=1
M302 271 267 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=12100 $Y=58500 $D=1
M303 272 38 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=12100 $Y=71850 $D=1
M304 273 94 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=12100 $Y=76300 $D=1
M305 274 39 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=12100 $Y=89650 $D=1
M306 275 95 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=12100 $Y=94100 $D=1
M307 450 90 268 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=12550 $Y=5100 $D=1
M308 451 91 269 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=12550 $Y=22900 $D=1
M309 452 92 270 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=12550 $Y=40700 $D=1
M310 453 93 271 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=12550 $Y=58500 $D=1
M311 GND! 94 450 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=13000 $Y=5100 $D=1
M312 GND! 95 451 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=13000 $Y=22900 $D=1
M313 GND! 96 452 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=13000 $Y=40700 $D=1
M314 GND! 89 453 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=13000 $Y=58500 $D=1
M315 97 272 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=13100 $Y=71850 $D=1
M316 102 273 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=13100 $Y=76300 $D=1
M317 98 274 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=13100 $Y=89650 $D=1
M318 103 275 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=13100 $Y=94100 $D=1
M319 108 268 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=13900 $Y=5100 $D=1
M320 99 269 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=13900 $Y=22900 $D=1
M321 100 270 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=13900 $Y=40700 $D=1
M322 101 271 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=13900 $Y=58500 $D=1
M323 280 213 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=14900 $Y=14000 $D=1
M324 281 35 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=14900 $Y=18450 $D=1
M325 282 99 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=14900 $Y=22900 $D=1
M326 283 214 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=14900 $Y=31800 $D=1
M327 284 36 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=14900 $Y=36250 $D=1
M328 285 100 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=14900 $Y=40700 $D=1
M329 286 215 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=14900 $Y=49600 $D=1
M330 287 37 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=14900 $Y=54050 $D=1
M331 288 101 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=14900 $Y=58500 $D=1
M332 289 216 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=14900 $Y=67400 $D=1
M333 290 217 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=14900 $Y=85200 $D=1
M334 291 218 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=14900 $Y=103000 $D=1
M335 292 219 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=14900 $Y=120800 $D=1
M336 454 57 280 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=15350 $Y=14000 $D=1
M337 455 58 283 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=15350 $Y=31800 $D=1
M338 456 59 286 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=15350 $Y=49600 $D=1
M339 457 60 289 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=15350 $Y=67400 $D=1
M340 458 61 290 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=15350 $Y=85200 $D=1
M341 459 62 291 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=15350 $Y=103000 $D=1
M342 460 63 292 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=15350 $Y=120800 $D=1
M343 GND! 99 454 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=15800 $Y=14000 $D=1
M344 GND! 100 455 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=15800 $Y=31800 $D=1
M345 GND! 101 456 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=15800 $Y=49600 $D=1
M346 GND! 102 457 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=15800 $Y=67400 $D=1
M347 GND! 103 458 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=15800 $Y=85200 $D=1
M348 GND! 96 459 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=15800 $Y=103000 $D=1
M349 GND! 89 460 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=15800 $Y=120800 $D=1
M350 104 281 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=15900 $Y=18450 $D=1
M351 110 282 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=15900 $Y=22900 $D=1
M352 105 284 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=15900 $Y=36250 $D=1
M353 112 285 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=15900 $Y=40700 $D=1
M354 106 287 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=15900 $Y=54050 $D=1
M355 114 288 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=15900 $Y=58500 $D=1
M356 109 280 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=16700 $Y=14000 $D=1
M357 111 283 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=16700 $Y=31800 $D=1
M358 113 286 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=16700 $Y=49600 $D=1
M359 115 289 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=16700 $Y=67400 $D=1
M360 116 290 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=16700 $Y=85200 $D=1
M361 117 291 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=16700 $Y=103000 $D=1
M362 118 292 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=16700 $Y=120800 $D=1
M363 300 151 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=-3800 $D=1
M364 301 108 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=5100 $D=1
M365 302 109 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=14000 $D=1
M366 303 110 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=22900 $D=1
M367 304 111 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=31800 $D=1
M368 305 112 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=40700 $D=1
M369 306 113 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=49600 $D=1
M370 307 114 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=58500 $D=1
M371 308 115 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=67400 $D=1
M372 309 102 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=76300 $D=1
M373 310 116 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=85200 $D=1
M374 311 103 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=94100 $D=1
M375 312 117 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=103000 $D=1
M376 313 96 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=111900 $D=1
M377 314 118 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=120800 $D=1
M378 315 89 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=17700 $Y=129700 $D=1
M379 461 41 300 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=18150 $Y=-3800 $D=1
M380 GND! 41 301 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=5100 $D=1
M381 GND! 33 302 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=14000 $D=1
M382 GND! 57 303 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=22900 $D=1
M383 GND! 104 304 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=31800 $D=1
M384 GND! 58 305 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=40700 $D=1
M385 GND! 105 306 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=49600 $D=1
M386 GND! 59 307 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=58500 $D=1
M387 GND! 106 308 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=67400 $D=1
M388 GND! 60 309 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=76300 $D=1
M389 GND! 97 310 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=85200 $D=1
M390 GND! 61 311 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=94100 $D=1
M391 GND! 98 312 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=103000 $D=1
M392 GND! 62 313 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=111900 $D=1
M393 GND! 107 314 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=120800 $D=1
M394 GND! 63 315 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=18150 $Y=129700 $D=1
M395 GND! 108 461 GND! NMOS_VTL L=5e-08 W=1e-07 AD=4e-14 AS=1.75e-14 PD=1e-06 PS=5.5e-07 $X=18600 $Y=-3800 $D=1
M396 GND! 301 S_15 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=5100 $D=1
M397 GND! 302 S_14 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=14000 $D=1
M398 GND! 303 S_13 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=22900 $D=1
M399 GND! 304 S_12 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=31800 $D=1
M400 GND! 305 S_11 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=40700 $D=1
M401 GND! 306 S_10 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=49600 $D=1
M402 GND! 307 S_9 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=58500 $D=1
M403 GND! 308 S_8 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=67400 $D=1
M404 GND! 309 S_7 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=76300 $D=1
M405 GND! 310 S_6 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=85200 $D=1
M406 GND! 311 S_5 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=94100 $D=1
M407 GND! 312 S_4 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=103000 $D=1
M408 GND! 313 S_3 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=111900 $D=1
M409 GND! 314 S_2 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=120800 $D=1
M410 GND! 315 S_1 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.5e-14 PD=5.5e-07 PS=5e-07 $X=19050 $Y=129700 $D=1
M411 Cout 300 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=4e-14 PD=5e-07 PS=1e-06 $X=19500 $Y=-3800 $D=1
M412 462 108 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=5100 $D=1
M413 463 109 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=14000 $D=1
M414 464 110 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=22900 $D=1
M415 465 111 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=31800 $D=1
M416 466 112 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=40700 $D=1
M417 467 113 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=49600 $D=1
M418 468 114 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=58500 $D=1
M419 469 115 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=67400 $D=1
M420 470 102 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=76300 $D=1
M421 471 116 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=85200 $D=1
M422 472 103 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=94100 $D=1
M423 473 117 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=103000 $D=1
M424 474 96 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=111900 $D=1
M425 475 118 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=120800 $D=1
M426 476 89 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.75e-14 AS=1.75e-14 PD=5.5e-07 PS=5.5e-07 $X=19500 $Y=129700 $D=1
M427 S_15 41 462 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=5100 $D=1
M428 S_14 33 463 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=14000 $D=1
M429 S_13 57 464 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=22900 $D=1
M430 S_12 104 465 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=31800 $D=1
M431 S_11 58 466 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=40700 $D=1
M432 S_10 105 467 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=49600 $D=1
M433 S_9 59 468 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=58500 $D=1
M434 S_8 106 469 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=67400 $D=1
M435 S_7 60 470 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=76300 $D=1
M436 S_6 97 471 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=85200 $D=1
M437 S_5 61 472 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=94100 $D=1
M438 S_4 98 473 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=103000 $D=1
M439 S_3 62 474 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=111900 $D=1
M440 S_2 107 475 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=120800 $D=1
M441 S_1 63 476 GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.75e-14 PD=5e-07 PS=5.5e-07 $X=19950 $Y=129700 $D=1
M442 349 A_15 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=-6950 $D=0
M443 120 A_15 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=-2500 $D=0
M444 350 A_14 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=1950 $D=0
M445 122 A_14 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=6400 $D=0
M446 351 A_13 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=10850 $D=0
M447 124 A_13 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=15300 $D=0
M448 352 A_12 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=19750 $D=0
M449 126 A_12 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=24200 $D=0
M450 353 A_11 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=28650 $D=0
M451 128 A_11 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=33100 $D=0
M452 354 A_10 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=37550 $D=0
M453 130 A_10 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=42000 $D=0
M454 355 A_9 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=46450 $D=0
M455 132 A_9 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=50900 $D=0
M456 356 A_8 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=55350 $D=0
M457 134 A_8 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=59800 $D=0
M458 357 A_7 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=64250 $D=0
M459 136 A_7 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=68700 $D=0
M460 358 A_6 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=73150 $D=0
M461 138 A_6 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=77600 $D=0
M462 359 A_5 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=82050 $D=0
M463 140 A_5 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=86500 $D=0
M464 360 A_4 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=90950 $D=0
M465 142 A_4 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=95400 $D=0
M466 361 A_3 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=99850 $D=0
M467 144 A_3 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=104300 $D=0
M468 362 A_2 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=108750 $D=0
M469 146 A_2 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=113200 $D=0
M470 363 A_1 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=117650 $D=0
M471 148 A_1 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=122100 $D=0
M472 364 A_0 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=126550 $D=0
M473 150 A_0 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=450 $Y=131000 $D=0
M474 119 B_15 349 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=-6950 $D=0
M475 VDD! B_15 120 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=-2500 $D=0
M476 121 B_14 350 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=1950 $D=0
M477 VDD! B_14 122 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=6400 $D=0
M478 123 B_13 351 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=10850 $D=0
M479 VDD! B_13 124 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=15300 $D=0
M480 125 B_12 352 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=19750 $D=0
M481 VDD! B_12 126 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=24200 $D=0
M482 127 B_11 353 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=28650 $D=0
M483 VDD! B_11 128 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=33100 $D=0
M484 129 B_10 354 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=37550 $D=0
M485 VDD! B_10 130 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=42000 $D=0
M486 131 B_9 355 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=46450 $D=0
M487 VDD! B_9 132 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=50900 $D=0
M488 133 B_8 356 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=55350 $D=0
M489 VDD! B_8 134 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=59800 $D=0
M490 135 B_7 357 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=64250 $D=0
M491 VDD! B_7 136 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=68700 $D=0
M492 137 B_6 358 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=73150 $D=0
M493 VDD! B_6 138 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=77600 $D=0
M494 139 B_5 359 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=82050 $D=0
M495 VDD! B_5 140 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=86500 $D=0
M496 141 B_4 360 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=90950 $D=0
M497 VDD! B_4 142 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=95400 $D=0
M498 143 B_3 361 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=99850 $D=0
M499 VDD! B_3 144 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=104300 $D=0
M500 145 B_2 362 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=108750 $D=0
M501 VDD! B_2 146 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=113200 $D=0
M502 147 B_1 363 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=117650 $D=0
M503 VDD! B_1 148 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=122100 $D=0
M504 149 B_0 364 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=126550 $D=0
M505 VDD! B_0 150 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=900 $Y=131000 $D=0
M506 160 119 41 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=-6950 $D=0
M507 161 121 33 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=1950 $D=0
M508 162 123 34 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=10850 $D=0
M509 163 125 35 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=19750 $D=0
M510 164 127 42 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=28650 $D=0
M511 165 129 36 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=37550 $D=0
M512 166 131 43 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=46450 $D=0
M513 167 133 37 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=55350 $D=0
M514 168 135 44 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=64250 $D=0
M515 169 137 38 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=73150 $D=0
M516 170 139 45 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=82050 $D=0
M517 171 141 39 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=90950 $D=0
M518 172 143 46 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=99850 $D=0
M519 173 145 40 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=108750 $D=0
M520 174 147 47 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=117650 $D=0
M521 175 149 55 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=1800 $Y=126550 $D=0
M522 151 120 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=-2500 $D=0
M523 152 122 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=6400 $D=0
M524 48 124 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=15300 $D=0
M525 153 126 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=24200 $D=0
M526 49 128 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=33100 $D=0
M527 154 130 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=42000 $D=0
M528 50 132 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=50900 $D=0
M529 155 134 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=59800 $D=0
M530 51 136 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=68700 $D=0
M531 156 138 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=77600 $D=0
M532 52 140 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=86500 $D=0
M533 157 142 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=95400 $D=0
M534 53 144 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=104300 $D=0
M535 158 146 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=113200 $D=0
M536 54 148 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=122100 $D=0
M537 159 150 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1900 $Y=131000 $D=0
M538 VDD! A_15 160 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=-6950 $D=0
M539 VDD! A_14 161 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=1950 $D=0
M540 VDD! A_13 162 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=10850 $D=0
M541 VDD! A_12 163 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=19750 $D=0
M542 VDD! A_11 164 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=28650 $D=0
M543 VDD! A_10 165 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=37550 $D=0
M544 VDD! A_9 166 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=46450 $D=0
M545 VDD! A_8 167 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=55350 $D=0
M546 VDD! A_7 168 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=64250 $D=0
M547 VDD! A_6 169 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=73150 $D=0
M548 VDD! A_5 170 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=82050 $D=0
M549 VDD! A_4 171 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=90950 $D=0
M550 VDD! A_3 172 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=99850 $D=0
M551 VDD! A_2 173 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=108750 $D=0
M552 VDD! A_1 174 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=117650 $D=0
M553 VDD! A_0 175 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=2250 $Y=126550 $D=0
M554 160 B_15 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=-6950 $D=0
M555 161 B_14 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=1950 $D=0
M556 162 B_13 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=10850 $D=0
M557 163 B_12 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=19750 $D=0
M558 164 B_11 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=28650 $D=0
M559 165 B_10 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=37550 $D=0
M560 166 B_9 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=46450 $D=0
M561 167 B_8 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=55350 $D=0
M562 168 B_7 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=64250 $D=0
M563 169 B_6 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=73150 $D=0
M564 170 B_5 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=82050 $D=0
M565 171 B_4 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=90950 $D=0
M566 172 B_3 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=99850 $D=0
M567 173 B_2 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=108750 $D=0
M568 174 B_1 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=117650 $D=0
M569 175 B_0 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=2700 $Y=126550 $D=0
M570 198 34 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=1950 $D=0
M571 205 152 176 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=6400 $D=0
M572 177 34 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=10850 $D=0
M573 178 48 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=15300 $D=0
M574 199 42 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=19750 $D=0
M575 206 153 179 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=24200 $D=0
M576 180 42 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=28650 $D=0
M577 181 49 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=33100 $D=0
M578 200 43 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=37550 $D=0
M579 207 154 182 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=42000 $D=0
M580 183 43 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=46450 $D=0
M581 184 50 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=50900 $D=0
M582 201 44 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=55350 $D=0
M583 208 155 185 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=59800 $D=0
M584 186 44 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=64250 $D=0
M585 187 51 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=68700 $D=0
M586 202 45 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=73150 $D=0
M587 209 156 188 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=77600 $D=0
M588 189 45 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=82050 $D=0
M589 190 52 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=86500 $D=0
M590 203 46 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=90950 $D=0
M591 210 157 191 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=95400 $D=0
M592 192 46 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=99850 $D=0
M593 193 53 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=104300 $D=0
M594 204 47 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=108750 $D=0
M595 211 158 194 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=113200 $D=0
M596 195 47 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=117650 $D=0
M597 196 54 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=3700 $Y=122100 $D=0
M598 212 159 197 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=3700 $Y=131000 $D=0
M599 VDD! 33 198 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4150 $Y=1950 $D=0
M600 VDD! 33 205 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=4150 $Y=6400 $D=0
M601 VDD! 35 199 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4150 $Y=19750 $D=0
M602 VDD! 35 206 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=4150 $Y=24200 $D=0
M603 VDD! 36 200 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4150 $Y=37550 $D=0
M604 VDD! 36 207 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=4150 $Y=42000 $D=0
M605 VDD! 37 201 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4150 $Y=55350 $D=0
M606 VDD! 37 208 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=4150 $Y=59800 $D=0
M607 VDD! 38 202 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4150 $Y=73150 $D=0
M608 VDD! 38 209 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=4150 $Y=77600 $D=0
M609 VDD! 39 203 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4150 $Y=90950 $D=0
M610 VDD! 39 210 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=4150 $Y=95400 $D=0
M611 VDD! 40 204 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4150 $Y=108750 $D=0
M612 VDD! 40 211 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=4150 $Y=113200 $D=0
M613 VDD! 55 212 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=4150 $Y=131000 $D=0
M614 205 48 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4600 $Y=6400 $D=0
M615 206 49 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4600 $Y=24200 $D=0
M616 207 50 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4600 $Y=42000 $D=0
M617 208 51 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4600 $Y=59800 $D=0
M618 209 52 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4600 $Y=77600 $D=0
M619 210 53 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4600 $Y=95400 $D=0
M620 211 54 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4600 $Y=113200 $D=0
M621 212 GND! VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=4600 $Y=131000 $D=0
M622 57 177 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=10850 $D=0
M623 213 178 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=15300 $D=0
M624 58 180 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=28650 $D=0
M625 214 181 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=33100 $D=0
M626 59 183 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=46450 $D=0
M627 215 184 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=50900 $D=0
M628 60 186 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=64250 $D=0
M629 216 187 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=68700 $D=0
M630 61 189 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=82050 $D=0
M631 217 190 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=86500 $D=0
M632 62 192 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=99850 $D=0
M633 218 193 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=104300 $D=0
M634 63 195 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=117650 $D=0
M635 219 196 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=4700 $Y=122100 $D=0
M636 64 198 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5150 $Y=1950 $D=0
M637 65 199 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5150 $Y=19750 $D=0
M638 66 200 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5150 $Y=37550 $D=0
M639 67 201 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5150 $Y=55350 $D=0
M640 68 202 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5150 $Y=73150 $D=0
M641 69 203 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5150 $Y=90950 $D=0
M642 70 204 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5150 $Y=108750 $D=0
M643 220 176 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5500 $Y=6400 $D=0
M644 71 179 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5500 $Y=24200 $D=0
M645 72 182 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5500 $Y=42000 $D=0
M646 73 185 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5500 $Y=59800 $D=0
M647 74 188 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5500 $Y=77600 $D=0
M648 75 191 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5500 $Y=95400 $D=0
M649 76 194 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5500 $Y=113200 $D=0
M650 77 197 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=5500 $Y=131000 $D=0
M651 230 65 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=1950 $D=0
M652 236 220 221 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=6400 $D=0
M653 231 66 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=19750 $D=0
M654 237 71 222 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=24200 $D=0
M655 232 67 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=37550 $D=0
M656 238 72 223 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=42000 $D=0
M657 233 68 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=55350 $D=0
M658 239 73 224 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=59800 $D=0
M659 234 69 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=73150 $D=0
M660 240 74 225 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=77600 $D=0
M661 235 70 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=90950 $D=0
M662 241 75 226 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=95400 $D=0
M663 242 76 227 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=6500 $Y=113200 $D=0
M664 228 55 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=6500 $Y=126550 $D=0
M665 229 77 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=6500 $Y=131000 $D=0
M666 VDD! 64 230 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=6950 $Y=1950 $D=0
M667 VDD! 64 236 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=6950 $Y=6400 $D=0
M668 VDD! 65 231 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=6950 $Y=19750 $D=0
M669 VDD! 65 237 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=6950 $Y=24200 $D=0
M670 VDD! 66 232 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=6950 $Y=37550 $D=0
M671 VDD! 66 238 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=6950 $Y=42000 $D=0
M672 VDD! 67 233 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=6950 $Y=55350 $D=0
M673 VDD! 67 239 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=6950 $Y=59800 $D=0
M674 VDD! 68 234 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=6950 $Y=73150 $D=0
M675 VDD! 68 240 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=6950 $Y=77600 $D=0
M676 VDD! 69 235 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=6950 $Y=90950 $D=0
M677 VDD! 69 241 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=6950 $Y=95400 $D=0
M678 VDD! 70 242 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=6950 $Y=113200 $D=0
M679 236 71 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=7400 $Y=6400 $D=0
M680 237 72 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=7400 $Y=24200 $D=0
M681 238 73 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=7400 $Y=42000 $D=0
M682 239 74 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=7400 $Y=59800 $D=0
M683 240 75 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=7400 $Y=77600 $D=0
M684 241 76 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=7400 $Y=95400 $D=0
M685 242 77 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=7400 $Y=113200 $D=0
M686 S_0 228 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=7500 $Y=126550 $D=0
M687 89 229 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=7500 $Y=131000 $D=0
M688 78 230 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=7950 $Y=1950 $D=0
M689 79 231 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=7950 $Y=19750 $D=0
M690 80 232 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=7950 $Y=37550 $D=0
M691 81 233 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=7950 $Y=55350 $D=0
M692 82 234 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=7950 $Y=73150 $D=0
M693 83 235 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=7950 $Y=90950 $D=0
M694 244 221 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=8300 $Y=6400 $D=0
M695 245 222 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=8300 $Y=24200 $D=0
M696 87 223 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=8300 $Y=42000 $D=0
M697 85 224 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=8300 $Y=59800 $D=0
M698 84 225 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=8300 $Y=77600 $D=0
M699 88 226 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=8300 $Y=95400 $D=0
M700 86 227 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=8300 $Y=113200 $D=0
M701 254 80 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=1950 $D=0
M702 258 244 246 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=6400 $D=0
M703 255 81 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=19750 $D=0
M704 259 245 247 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=24200 $D=0
M705 256 82 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=37550 $D=0
M706 260 87 248 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=42000 $D=0
M707 257 83 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=55350 $D=0
M708 261 85 249 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=59800 $D=0
M709 262 84 250 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=77600 $D=0
M710 263 88 251 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=9300 $Y=95400 $D=0
M711 252 40 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=9300 $Y=108750 $D=0
M712 253 86 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=9300 $Y=113200 $D=0
M713 VDD! 78 254 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=9750 $Y=1950 $D=0
M714 VDD! 78 258 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=9750 $Y=6400 $D=0
M715 VDD! 79 255 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=9750 $Y=19750 $D=0
M716 VDD! 79 259 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=9750 $Y=24200 $D=0
M717 VDD! 80 256 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=9750 $Y=37550 $D=0
M718 VDD! 80 260 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=9750 $Y=42000 $D=0
M719 VDD! 81 257 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=9750 $Y=55350 $D=0
M720 VDD! 81 261 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=9750 $Y=59800 $D=0
M721 VDD! 82 262 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=9750 $Y=77600 $D=0
M722 VDD! 83 263 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=9750 $Y=95400 $D=0
M723 258 87 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=10200 $Y=6400 $D=0
M724 259 85 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=10200 $Y=24200 $D=0
M725 260 84 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=10200 $Y=42000 $D=0
M726 261 88 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=10200 $Y=59800 $D=0
M727 262 86 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=10200 $Y=77600 $D=0
M728 263 89 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=10200 $Y=95400 $D=0
M729 107 252 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=10300 $Y=108750 $D=0
M730 96 253 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=10300 $Y=113200 $D=0
M731 90 254 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=10750 $Y=1950 $D=0
M732 91 255 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=10750 $Y=19750 $D=0
M733 92 256 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=10750 $Y=37550 $D=0
M734 93 257 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=10750 $Y=55350 $D=0
M735 264 246 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=11100 $Y=6400 $D=0
M736 265 247 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=11100 $Y=24200 $D=0
M737 266 248 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=11100 $Y=42000 $D=0
M738 267 249 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=11100 $Y=59800 $D=0
M739 94 250 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=11100 $Y=77600 $D=0
M740 95 251 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=11100 $Y=95400 $D=0
M741 276 264 268 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=12100 $Y=6400 $D=0
M742 277 265 269 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=12100 $Y=24200 $D=0
M743 278 266 270 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=12100 $Y=42000 $D=0
M744 279 267 271 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=12100 $Y=59800 $D=0
M745 272 38 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=12100 $Y=73150 $D=0
M746 273 94 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=12100 $Y=77600 $D=0
M747 274 39 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=12100 $Y=90950 $D=0
M748 275 95 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=12100 $Y=95400 $D=0
M749 VDD! 90 276 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=12550 $Y=6400 $D=0
M750 VDD! 91 277 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=12550 $Y=24200 $D=0
M751 VDD! 92 278 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=12550 $Y=42000 $D=0
M752 VDD! 93 279 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=12550 $Y=59800 $D=0
M753 276 94 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=13000 $Y=6400 $D=0
M754 277 95 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=13000 $Y=24200 $D=0
M755 278 96 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=13000 $Y=42000 $D=0
M756 279 89 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=13000 $Y=59800 $D=0
M757 97 272 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=13100 $Y=73150 $D=0
M758 102 273 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=13100 $Y=77600 $D=0
M759 98 274 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=13100 $Y=90950 $D=0
M760 103 275 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=13100 $Y=95400 $D=0
M761 108 268 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=13900 $Y=6400 $D=0
M762 99 269 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=13900 $Y=24200 $D=0
M763 100 270 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=13900 $Y=42000 $D=0
M764 101 271 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=13900 $Y=59800 $D=0
M765 293 213 280 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=14900 $Y=15300 $D=0
M766 281 35 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=14900 $Y=19750 $D=0
M767 282 99 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=14900 $Y=24200 $D=0
M768 294 214 283 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=14900 $Y=33100 $D=0
M769 284 36 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=14900 $Y=37550 $D=0
M770 285 100 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=14900 $Y=42000 $D=0
M771 295 215 286 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=14900 $Y=50900 $D=0
M772 287 37 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=14900 $Y=55350 $D=0
M773 288 101 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=14900 $Y=59800 $D=0
M774 296 216 289 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=14900 $Y=68700 $D=0
M775 297 217 290 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=14900 $Y=86500 $D=0
M776 298 218 291 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=14900 $Y=104300 $D=0
M777 299 219 292 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=14900 $Y=122100 $D=0
M778 VDD! 57 293 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=15350 $Y=15300 $D=0
M779 VDD! 58 294 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=15350 $Y=33100 $D=0
M780 VDD! 59 295 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=15350 $Y=50900 $D=0
M781 VDD! 60 296 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=15350 $Y=68700 $D=0
M782 VDD! 61 297 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=15350 $Y=86500 $D=0
M783 VDD! 62 298 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=15350 $Y=104300 $D=0
M784 VDD! 63 299 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=15350 $Y=122100 $D=0
M785 293 99 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=15800 $Y=15300 $D=0
M786 294 100 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=15800 $Y=33100 $D=0
M787 295 101 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=15800 $Y=50900 $D=0
M788 296 102 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=15800 $Y=68700 $D=0
M789 297 103 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=15800 $Y=86500 $D=0
M790 298 96 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=15800 $Y=104300 $D=0
M791 299 89 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=15800 $Y=122100 $D=0
M792 104 281 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=15900 $Y=19750 $D=0
M793 110 282 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=15900 $Y=24200 $D=0
M794 105 284 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=15900 $Y=37550 $D=0
M795 112 285 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=15900 $Y=42000 $D=0
M796 106 287 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=15900 $Y=55350 $D=0
M797 114 288 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=15900 $Y=59800 $D=0
M798 109 280 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=16700 $Y=15300 $D=0
M799 111 283 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=16700 $Y=33100 $D=0
M800 113 286 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=16700 $Y=50900 $D=0
M801 115 289 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=16700 $Y=68700 $D=0
M802 116 290 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=16700 $Y=86500 $D=0
M803 117 291 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=16700 $Y=104300 $D=0
M804 118 292 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=16700 $Y=122100 $D=0
M805 316 151 300 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=-2500 $D=0
M806 365 108 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=6400 $D=0
M807 366 109 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=15300 $D=0
M808 367 110 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=24200 $D=0
M809 368 111 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=33100 $D=0
M810 369 112 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=42000 $D=0
M811 370 113 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=50900 $D=0
M812 371 114 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=59800 $D=0
M813 372 115 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=68700 $D=0
M814 373 102 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=77600 $D=0
M815 374 116 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=86500 $D=0
M816 375 103 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=95400 $D=0
M817 376 117 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=104300 $D=0
M818 377 96 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=113200 $D=0
M819 378 118 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=122100 $D=0
M820 379 89 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=17700 $Y=131000 $D=0
M821 VDD! 41 316 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=18150 $Y=-2500 $D=0
M822 301 41 365 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=6400 $D=0
M823 302 33 366 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=15300 $D=0
M824 303 57 367 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=24200 $D=0
M825 304 104 368 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=33100 $D=0
M826 305 58 369 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=42000 $D=0
M827 306 105 370 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=50900 $D=0
M828 307 59 371 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=59800 $D=0
M829 308 106 372 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=68700 $D=0
M830 309 60 373 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=77600 $D=0
M831 310 97 374 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=86500 $D=0
M832 311 61 375 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=95400 $D=0
M833 312 98 376 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=104300 $D=0
M834 313 62 377 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=113200 $D=0
M835 314 107 378 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=122100 $D=0
M836 315 63 379 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18150 $Y=131000 $D=0
M837 316 108 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=18600 $Y=-2500 $D=0
M838 320 301 S_15 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=6400 $D=0
M839 322 302 S_14 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=15300 $D=0
M840 324 303 S_13 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=24200 $D=0
M841 326 304 S_12 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=33100 $D=0
M842 328 305 S_11 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=42000 $D=0
M843 330 306 S_10 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=50900 $D=0
M844 332 307 S_9 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=59800 $D=0
M845 334 308 S_8 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=68700 $D=0
M846 336 309 S_7 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=77600 $D=0
M847 338 310 S_6 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=86500 $D=0
M848 340 311 S_5 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=95400 $D=0
M849 342 312 S_4 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=104300 $D=0
M850 344 313 S_3 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=113200 $D=0
M851 346 314 S_2 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=122100 $D=0
M852 348 315 S_1 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3e-14 PD=7.5e-07 PS=7e-07 $X=19050 $Y=131000 $D=0
M853 Cout 300 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=19500 $Y=-2500 $D=0
M854 VDD! 108 320 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=6400 $D=0
M855 VDD! 109 322 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=15300 $D=0
M856 VDD! 110 324 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=24200 $D=0
M857 VDD! 111 326 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=33100 $D=0
M858 VDD! 112 328 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=42000 $D=0
M859 VDD! 113 330 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=50900 $D=0
M860 VDD! 114 332 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=59800 $D=0
M861 VDD! 115 334 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=68700 $D=0
M862 VDD! 102 336 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=77600 $D=0
M863 VDD! 116 338 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=86500 $D=0
M864 VDD! 103 340 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=95400 $D=0
M865 VDD! 117 342 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=104300 $D=0
M866 VDD! 96 344 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=113200 $D=0
M867 VDD! 118 346 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=122100 $D=0
M868 VDD! 89 348 VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3.5e-14 AS=3.5e-14 PD=7.5e-07 PS=7.5e-07 $X=19500 $Y=131000 $D=0
M869 320 41 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=6400 $D=0
M870 322 33 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=15300 $D=0
M871 324 57 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=24200 $D=0
M872 326 104 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=33100 $D=0
M873 328 58 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=42000 $D=0
M874 330 105 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=50900 $D=0
M875 332 59 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=59800 $D=0
M876 334 106 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=68700 $D=0
M877 336 60 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=77600 $D=0
M878 338 97 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=86500 $D=0
M879 340 61 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=95400 $D=0
M880 342 98 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=104300 $D=0
M881 344 62 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=113200 $D=0
M882 346 107 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=122100 $D=0
M883 348 63 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3.5e-14 PD=7e-07 PS=7.5e-07 $X=19950 $Y=131000 $D=0
.ENDS
***************************************
