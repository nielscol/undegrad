`timescale 1ns / 1ps
module divider(one_hz, clock);
	input clock;
	output one_hz;

	

endmodule
