A SIMPLE AC RUN
.OPTIONS LIST NODE POST
.TRAN 10U 10m
.PRINT TRAN V(1) V(2) I(R2)
V1 1 0 PULSE 0 1 0N 0N 20 10U 10U 
R1 1 2 1k
C1 2 0 1U
.END
