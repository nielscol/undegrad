A SIMPLE AC RUN
.OPTIONS LIST NODE POST
.AC DEC 10 10 100k
.PRINT AC V(1) V(2) I(R2)
V1 1 0 AC 1
R1 1 2 1k
C1 2 0 1U
.END
