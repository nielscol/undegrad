.GLOBAL VDD! 
   
C100 S_0 0 50E-15 M=1.0
C101 S_1 0 50E-15 M=1.0
C102 S_2 0 50E-15 M=1.0
C103 S_3 0 50E-15 M=1.0
C104 S_4 0 50E-15 M=1.0
C105 S_5 0 50E-15 M=1.0
C106 S_6 0 50E-15 M=1.0
C107 S_7 0 50E-15 M=1.0
C108 S_8 0 50E-15 M=1.0
C109 S_9 0 50E-15 M=1.0
C110 S_10 0 50E-15 M=1.0
C111 S_11 0 50E-15 M=1.0
C112 S_12 0 50E-15 M=1.0
C113 S_13 0 50E-15 M=1.0
C114 S_14 0 50E-15 M=1.0
C115 S_15 0 50E-15 M=1.0
C116 Cout 0 50E-15 M=1.0


XI170 A_BAR_0 A_BAR_1 A_BAR_2 A_BAR_3 A_BAR_4 A_BAR_5 A_BAR_6 A_BAR_7 A_BAR_8 A_BAR_9 A_BAR_10 A_BAR_11 A_BAR_12 A_BAR_13 A_BAR_14 A_BAR_15 
+AIN_0 AIN_1 AIN_2 AIN_3 AIN_4 AIN_5 AIN_6 AIN_7 AIN_8 AIN_9 AIN_10 AIN_11 AIN_12 AIN_13 AIN_14 AIN_15 INPUTBUF_G120 
XI180 A_0 A_1 A_2 A_3 A_4 A_5 A_6 A_7 A_8 A_9 A_10 A_11 A_12 A_13 A_14 A_15
+A_BAR_0 A_BAR_1 A_BAR_2 A_BAR_3 A_BAR_4 A_BAR_5 A_BAR_6 A_BAR_7 A_BAR_8 A_BAR_9 A_BAR_10 A_BAR_11 A_BAR_12 A_BAR_13 A_BAR_14 A_BAR_15 INPUTBUF_G120 

XI190 B_BAR_0 B_BAR_1 B_BAR_2 B_BAR_3 B_BAR_4 B_BAR_5 B_BAR_6 B_BAR_7 B_BAR_8 B_BAR_9 B_BAR_10 B_BAR_11 B_BAR_12 B_BAR_13 B_BAR_14 B_BAR_15 
+BIN_0 BIN_1 BIN_2 BIN_3 BIN_4 BIN_5 BIN_6 BIN_7 BIN_8 BIN_9 BIN_10 BIN_11 BIN_12 BIN_13 BIN_14 BIN_15 INPUTBUF_G120 
XI200 B_0 B_1 B_2 B_3 B_4 B_5 B_6 B_7 B_8 B_9 B_10 B_11 B_12 B_13 B_14 B_15
+B_BAR_0 B_BAR_1 B_BAR_2 B_BAR_3 B_BAR_4 B_BAR_5 B_BAR_6 B_BAR_7 B_BAR_8 B_BAR_9 B_BAR_10 B_BAR_11 B_BAR_12 B_BAR_13 B_BAR_14 B_BAR_15 INPUTBUF_G120 



.SUBCKT INV_G200 IN OUT 
m0 OUT IN 0 0 NMOS_VTL L=50e-9 W=200e-9
m2 OUT IN VDD! VDD! PMOS_VTL L=50e-9 W=300e-9
.ENDS INV_G200
 
.SUBCKT INPUTBUF_G120 OUT_0 OUT_1 OUT_2 OUT_3 OUT_4 OUT_5 OUT_6 OUT_7 OUT_8 OUT_9 OUT_10 OUT_11 OUT_12 OUT_13 OUT_14 OUT_15
+IN_0 IN_1 IN_2 IN_3 IN_4 IN_5 IN_6 IN_7 IN_8 IN_9 IN_10 IN_11 IN_12 IN_13 IN_14 IN_15 
XI15 IN_15 OUT_15 INV_G200 
XI14 IN_14 OUT_14 INV_G200 
XI13 IN_13 OUT_13 INV_G200 
XI12 IN_12 OUT_12 INV_G200 
XI11 IN_11 OUT_11 INV_G200 
XI10 IN_10 OUT_10 INV_G200 
XI9 IN_9 OUT_9 INV_G200 
XI8 IN_8 OUT_8 INV_G200 
XI7 IN_7 OUT_7 INV_G200 
XI6 IN_6 OUT_6 INV_G200 
XI5 IN_5 OUT_5 INV_G200 
XI4 IN_4 OUT_4 INV_G200 
XI3 IN_3 OUT_3 INV_G200 
XI2 IN_2 OUT_2 INV_G200 
XI1 IN_1 OUT_1 INV_G200 
XI0 IN_0 OUT_0 INV_G200 
.ENDS INPUTBUF_G120 

