* SPICE NETLIST
***************************************

.SUBCKT PG_buffer Pi Gi GND! VDD! Po Go
** N=8 EP=6 IP=0 FDC=8
M0 3 Pi GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=450 $Y=650 $D=1
M1 4 Gi GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=450 $Y=5100 $D=1
M2 Po 3 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1450 $Y=650 $D=1
M3 Go 4 GND! GND! NMOS_VTL L=5e-08 W=1e-07 AD=1.5e-14 AS=1.5e-14 PD=5e-07 PS=5e-07 $X=1450 $Y=5100 $D=1
M4 3 Pi VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=450 $Y=1950 $D=0
M5 4 Gi VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=450 $Y=6400 $D=0
M6 Po 3 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1450 $Y=1950 $D=0
M7 Go 4 VDD! VDD! PMOS_VTL L=5e-08 W=2e-07 AD=3e-14 AS=3e-14 PD=7e-07 PS=7e-07 $X=1450 $Y=6400 $D=0
.ENDS
***************************************
