*TEST 16-BIT ADDER
.TEMP 25
.OPTIONS ACCURATE
.OPTIONS POST=2
.OPTIONS MEASFORM=1

.INCLUDE '~/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/NMOS_VTL.inc'
.INCLUDE '~/FreePDK45/ncsu_basekit/models/hspice/tran_models/models_nom/PMOS_VTL.inc' 

.INCLUDE adder16b.sp
.INCLUDE testadder16b.sp
* YOU SHOULD CHECK DIFFERENT INPUT PATTERNS FOR
* MAXIMUM DELAY
.VEC 'digital_vector_delay'
.PARAM PERIOD = 4NS
.PARAM T0= 0.1NS
.PARAM T1= T0+PERIOD
.PARAM T2= T1+0.1NS
.PARAM STEP= 1PS

VDD   VDD! 0 1.1
VGND  GND! 0 0

.TRAN STEP T2

* YOU SHOULD MAKE SURE THAT YOU ARE MEASURING THE CORRECT SIGNAL FOR MAXIMUM DELAY. BELOW IS JUST AN EXAMPLE.
.MEASURE TRAN DELAY_MAX TRIG V(A_0) VAL= 0.55 RISE=1 TARG V(Cout) VAL= 0.55 RISE=1

.END








